module collision

import vector2

struct Collision {
	pos vector2.vector2
	rad f32
}

pub fn check() {
	
}
